`ifndef CONFIG_VH		// Guard prevents header file from being included more than once
`define CONFIG_VH

`define FEATURE_MULT
// `define FEATURE_DIV
// `define FEATURE_XILINX_DATAMEM_IP_GEN

`define REPO_LOCATION        "T:/Files/Projects/RV32IMC-Repo/pipelined-RV32IMC/"
`define TEST_LOCATION        "assembly-tests/riscv-compliance/"

`endif